module ROM(
    input clka,
    input [5:0] addra,
    output reg[31:0] douta
    );
    reg[31:0] ins_regs[0:63];
    initial begin
        ins_regs[0] = 32'b00000000000000000000100000100111;
        ins_regs[1] = 32'b00000000000000010001000000101011;
        ins_regs[2] = 32'b00000000010000100001100000100000;
        ins_regs[3] = 32'b00000000011000100010000000100000;
        ins_regs[4] = 32'b00000000100000110010100000100000;
        ins_regs[5] = 32'b00000000101000110011000000100000;
        ins_regs[6] = 32'b00000000010001100011100000000100;
        ins_regs[7] = 32'b00000000101001100100100000100000;
        ins_regs[8] = 32'b00000001001001100100000000000100;
        ins_regs[9] = 32'b00000000001010000100100000100110;
        ins_regs[10] = 32'b00000001001000010101000000100000;
        ins_regs[11] = 32'b00000001000001110101100000100010;
        ins_regs[12] = 32'b00000000111010000110000000100010;
        ins_regs[13] = 32'b00000001001011000110100000100100;
        ins_regs[14] = 32'b00000001001011000111000000100101;
    end
    always@(posedge clka) begin
        douta = ins_regs[addra];
    end
endmodule
